LIBRARY IEEE;
use IEEE.std_logic_1164.all;

entity part4 is
    port (
        D: in std_logic;
        Clk: in std_logic;
        Qb1: out std_logic;
        Qa1: out std_logic;
        Qb2: out std_logic;
        Qa2: out std_logic;
        Qb3: out std_logic;
        Qa3: out std_logic
    );
end entity part4;

architecture Behaviour of part4 is
begin   
    process(D, Clk)
    begin
        if Clk = '1' then
            Qb1 <= D;
            Qa1 <= not D;
        end if;
        if rising_edge(Clk) then
            Qb2 <= D;
            Qa2 <= not D;
        end if;
        if falling_edge(Clk) then
            Qb3 <= D;
            Qa3 <= not D;
        end if;
    end process;
end architecture;
